module love;

endmodule
