module love;
  $display("");
endmodule
